module conv_top_test #(
    parameter DATA_WIDTH = 16,    // Half-precision float width
    parameter KERNEL_SIZE = 5,
    parameter STRIDE = 1,
    parameter PADDING = 1,
    localparam DATA_ARRAY = DATA_WIDTH * KERNEL_SIZE,
    parameter CONV_OUTPUT = 16,   // Changed to match DATA_WIDTH for FP16
    parameter IMAGE_SIZE = 28     
)(
    input logic clk,
    input logic rst,

    // BRAM_PS Interface
    input logic [255:0] data_out,   
    output logic [11:0] bram_addr_a_ps,
    // output logic write_enable,
    // output logic bram_en_a_ps,


    input logic start,
    output logic done,
    // output logic done_1,
    // output logic done_2,
    // output logic done_3,
    output logic [DATA_WIDTH-1:0] data_out_0, // Output convolution result
    output logic [DATA_WIDTH-1:0] data_out_1,
    output logic [DATA_WIDTH-1:0] data_out_2,
    output logic [DATA_WIDTH-1:0] data_out_3,
    output logic [DATA_WIDTH-1:0] data_out_4,
    output logic [DATA_WIDTH-1:0] data_out_5,
    output logic [DATA_WIDTH-1:0] data_out_6,
    output logic [DATA_WIDTH-1:0] data_out_7,
    output logic [DATA_WIDTH-1:0] data_out_8,
    output logic [DATA_WIDTH-1:0] data_out_9,
    output logic [DATA_WIDTH-1:0] data_out_10,
    output logic [DATA_WIDTH-1:0] data_out_11,
    output logic [DATA_WIDTH-1:0] data_out_12,
    output logic [DATA_WIDTH-1:0] data_out_13,
    output logic [DATA_WIDTH-1:0] data_out_14,
    output logic [DATA_WIDTH-1:0] data_out_15,
    output logic [DATA_WIDTH-1:0] data_out_16,
    output logic [DATA_WIDTH-1:0] data_out_17,
    output logic [DATA_WIDTH-1:0] data_out_18,
    output logic [DATA_WIDTH-1:0] data_out_19,
    output logic [DATA_WIDTH-1:0] data_out_20,
    output logic [DATA_WIDTH-1:0] data_out_21,
    output logic [DATA_WIDTH-1:0] data_out_22,
    output logic [DATA_WIDTH-1:0] data_out_23,
    // output logic [DATA_WIDTH-1:0] data_out_24,
    // output logic [DATA_WIDTH-1:0] data_out_25,
    // output logic [DATA_WIDTH-1:0] data_out_26,
    // output logic [DATA_WIDTH-1:0] data_out_27,
    // output logic [DATA_WIDTH-1:0] data_out_28,
    // output logic [DATA_WIDTH-1:0] data_out_29,
    // output logic [DATA_WIDTH-1:0] data_out_30,
    // output logic [DATA_WIDTH-1:0] data_out_31,
    // output logic [DATA_WIDTH-1:0] data_out_32,
    // output logic [DATA_WIDTH-1:0] data_out_33,
    // output logic [DATA_WIDTH-1:0] data_out_34,
    // output logic [DATA_WIDTH-1:0] data_out_35,
    // output logic [DATA_WIDTH-1:0] data_out_36,
    // output logic [DATA_WIDTH-1:0] data_out_37,
    // output logic [DATA_WIDTH-1:0] data_out_38,
    // output logic [DATA_WIDTH-1:0] data_out_39,
    // output logic [DATA_WIDTH-1:0] data_out_40,
    // output logic [DATA_WIDTH-1:0] data_out_41,
    // output logic [DATA_WIDTH-1:0] data_out_42,
    // output logic [DATA_WIDTH-1:0] data_out_43,
    // output logic [DATA_WIDTH-1:0] data_out_44,
    // output logic [DATA_WIDTH-1:0] data_out_45,
    // output logic [DATA_WIDTH-1:0] data_out_46,
    // output logic [DATA_WIDTH-1:0] data_out_47,
    // output logic [DATA_WIDTH-1:0] data_out_48,
    // output logic [DATA_WIDTH-1:0] data_out_49,
    // output logic [DATA_WIDTH-1:0] data_out_50,
    // output logic [DATA_WIDTH-1:0] data_out_51,
    // output logic [DATA_WIDTH-1:0] data_out_52,
    // output logic [DATA_WIDTH-1:0] data_out_53,
    // output logic [DATA_WIDTH-1:0] data_out_54,
    // output logic [DATA_WIDTH-1:0] data_out_55,
    // output logic [DATA_WIDTH-1:0] data_out_56,
    // output logic [DATA_WIDTH-1:0] data_out_57,
    // output logic [DATA_WIDTH-1:0] data_out_58,
    // output logic [DATA_WIDTH-1:0] data_out_59,
    // output logic [DATA_WIDTH-1:0] data_out_60,
    // output logic [DATA_WIDTH-1:0] data_out_61,
    // output logic [DATA_WIDTH-1:0] data_out_62,
    // output logic [DATA_WIDTH-1:0] data_out_63,
    // output logic [DATA_WIDTH-1:0] data_out_64,
    // output logic [DATA_WIDTH-1:0] data_out_65,
    // output logic [DATA_WIDTH-1:0] data_out_66,
    // output logic [DATA_WIDTH-1:0] data_out_67,
    // output logic [DATA_WIDTH-1:0] data_out_68,
    // output logic [DATA_WIDTH-1:0] data_out_69,
    // output logic [DATA_WIDTH-1:0] data_out_70,
    // output logic [DATA_WIDTH-1:0] data_out_71,
    // output logic [DATA_WIDTH-1:0] data_out_72,
    // output logic [DATA_WIDTH-1:0] data_out_73,
    // output logic [DATA_WIDTH-1:0] data_out_74,
    // output logic [DATA_WIDTH-1:0] data_out_75,
    // output logic [DATA_WIDTH-1:0] data_out_76,
    // output logic [DATA_WIDTH-1:0] data_out_77,
    // output logic [DATA_WIDTH-1:0] data_out_78,
    // output logic [DATA_WIDTH-1:0] data_out_79,
    // output logic [DATA_WIDTH-1:0] data_out_80,
    // output logic [DATA_WIDTH-1:0] data_out_81,
    // output logic [DATA_WIDTH-1:0] data_out_82,
    // output logic [DATA_WIDTH-1:0] data_out_83,
    // output logic [DATA_WIDTH-1:0] data_out_84,
    // output logic [DATA_WIDTH-1:0] data_out_85,
    // output logic [DATA_WIDTH-1:0] data_out_86,
    // output logic [DATA_WIDTH-1:0] data_out_87,
    // output logic [DATA_WIDTH-1:0] data_out_88,
    // output logic [DATA_WIDTH-1:0] data_out_89,
    // output logic [DATA_WIDTH-1:0] data_out_90,
    // output logic [DATA_WIDTH-1:0] data_out_91,
    // output logic [DATA_WIDTH-1:0] data_out_92,
    // output logic [DATA_WIDTH-1:0] data_out_93,
    // output logic [DATA_WIDTH-1:0] data_out_94,
    // output logic [DATA_WIDTH-1:0] data_out_95,
    output logic valid_out,
    output logic keep_top
);


// assign bram_en_a_ps = 1'b1; // Read enable signal for BRAM
//logic [15:0] output_data [IMAGE_SIZE-KERNEL_SIZE:0];

edge_detection_test #(
    .DATA_WIDTH(DATA_WIDTH),
    .KERNEL_SIZE(KERNEL_SIZE),
    .STRIDE(STRIDE),
    .PADDING(PADDING),
    .CONV_OUTPUT(CONV_OUTPUT),
    .IMAGE_SIZE(IMAGE_SIZE)
) edge_detect (
    .clk(clk),
    .rst(rst),
    .start(start),
    .write_enable(), // Unconnected - not used
    .read_enable(),  // Unconnected - not used
    .data_in(data_out[255:0]), // Input image data
    .data_out_0(data_out_0), // Output convolution result
    .data_out_1(data_out_1),
    .data_out_2(data_out_2),
    .data_out_3(data_out_3),
    .data_out_4(data_out_4),
    .data_out_5(data_out_5),
    .data_out_6(data_out_6),
    .data_out_7(data_out_7),
    .data_out_8(data_out_8),
    .data_out_9(data_out_9),
    .data_out_10(data_out_10),
    .data_out_11(data_out_11),
    .data_out_12(data_out_12),
    .data_out_13(data_out_13),
    .data_out_14(data_out_14),
    .data_out_15(data_out_15),
    .data_out_16(data_out_16),
    .data_out_17(data_out_17),
    .data_out_18(data_out_18),
    .data_out_19(data_out_19),
    .data_out_20(data_out_20),
    .data_out_21(data_out_21),
    .data_out_22(data_out_22),
    .data_out_23(data_out_23),
    .addr(bram_addr_a_ps), // Address output
    .done(done),
    .valid_out_col(valid_out),
    .out_col_num(),  // Unconnected - not used

    .keep(keep_top)
);

// edge_detection #(
//     .DATA_WIDTH(DATA_WIDTH),
//     .KERNEL_SIZE(KERNEL_SIZE),
//     .STRIDE(STRIDE),
//     .PADDING(PADDING),
//     .CONV_OUTPUT(CONV_OUTPUT),
//     .IMAGE_SIZE(IMAGE_SIZE)
// ) edge_detect_1 (
//     .clk(clk),
//     .rst(rst),
//     .start(start),
//     // .write_enable(write_enable),
//     // .read_enable(read_enable),
//     .data_in(data_out[255:0]),
//     .data_out_0(data_out_24),
//     .data_out_1(data_out_25),
//     .data_out_2(data_out_26),
//     .data_out_3(data_out_27),
//     .data_out_4(data_out_28),
//     .data_out_5(data_out_29),
//     .data_out_6(data_out_30),
//     .data_out_7(data_out_31),
//     .data_out_8(data_out_32),
//     .data_out_9(data_out_33),
//     .data_out_10(data_out_34),
//     .data_out_11(data_out_35),
//     .data_out_12(data_out_36),
//     .data_out_13(data_out_37),
//     .data_out_14(data_out_38),
//     .data_out_15(data_out_39),
//     .data_out_16(data_out_40),
//     .data_out_17(data_out_41),
//     .data_out_18(data_out_42),
//     .data_out_19(data_out_43),
//     .data_out_20(data_out_44),
//     .data_out_21(data_out_45),
//     .data_out_22(data_out_46),
//     .data_out_23(data_out_47),
//     // .addr(), // Unconnected address
//     .done(done_1)
// //    .valid_in()
// );

// edge_detection #(
//     .DATA_WIDTH(DATA_WIDTH),
//     .KERNEL_SIZE(KERNEL_SIZE),
//     .STRIDE(STRIDE),
//     .PADDING(PADDING),
//     .CONV_OUTPUT(CONV_OUTPUT),
//     .IMAGE_SIZE(IMAGE_SIZE)
// ) edge_detect_2 (
//     .clk(clk),
//     .rst(rst),
//     .start(start),
//     // .write_enable(write_enable),
//     // .read_enable(read_enable),
//     .data_in(data_out[255:0]),
//     .data_out_0(data_out_48),
//     .data_out_1(data_out_49),
//     .data_out_2(data_out_50),
//     .data_out_3(data_out_51),
//     .data_out_4(data_out_52),
//     .data_out_5(data_out_53),
//     .data_out_6(data_out_54),
//     .data_out_7(data_out_55),
//     .data_out_8(data_out_56),
//     .data_out_9(data_out_57),
//     .data_out_10(data_out_58),
//     .data_out_11(data_out_59),
//     .data_out_12(data_out_60),
//     .data_out_13(data_out_61),
//     .data_out_14(data_out_62),
//     .data_out_15(data_out_63),
//     .data_out_16(data_out_64),
//     .data_out_17(data_out_65),
//     .data_out_18(data_out_66),
//     .data_out_19(data_out_67),
//     .data_out_20(data_out_68),
//     .data_out_21(data_out_69),
//     .data_out_22(data_out_70),
//     .data_out_23(data_out_71),
//     // .addr(),
//     .done(done_2)
// //    .valid_out_col()
// );

// edge_detection #(
//     .DATA_WIDTH(DATA_WIDTH),
//     .KERNEL_SIZE(KERNEL_SIZE),
//     .STRIDE(STRIDE),
//     .PADDING(PADDING),
//     .CONV_OUTPUT(CONV_OUTPUT),
//     .IMAGE_SIZE(IMAGE_SIZE)
// ) edge_detect_3 (
//     .clk(clk),
//     .rst(rst),
//     .start(start),
//     // .write_enable(write_enable),
//     // .read_enable(read_enable),
//     .data_in(data_out[255:0]),
//     .data_out_0(data_out_72),
//     .data_out_1(data_out_73),
//     .data_out_2(data_out_74),
//     .data_out_3(data_out_75),
//     .data_out_4(data_out_76),
//     .data_out_5(data_out_77),
//     .data_out_6(data_out_78),
//     .data_out_7(data_out_79),
//     .data_out_8(data_out_80),
//     .data_out_9(data_out_81),
//     .data_out_10(data_out_82),
//     .data_out_11(data_out_83),
//     .data_out_12(data_out_84),
//     .data_out_13(data_out_85),
//     .data_out_14(data_out_86),
//     .data_out_15(data_out_87),
//     .data_out_16(data_out_88),
//     .data_out_17(data_out_89),
//     .data_out_18(data_out_90),
//     .data_out_19(data_out_91),
//     .data_out_20(data_out_92),
//     .data_out_21(data_out_93),
//     .data_out_22(data_out_94),
//     .data_out_23(data_out_95),
//     // .addr(),
//     .done(done_3)
// //    .valid_in()
// );



// bram #() bram_inst (
//     .clk(clk),
//     .address(addr),
//     .write_enable(write_enable), // Assuming write_enable is controlled by start signal
//     .read_enable(read_enable), // Read when not writing
//     .data_in(data_in),
//     .data_out(data_out)
// );

endmodule

// Convolutional Layer Parameters

localparam [15:0] KERNELS[0:3][0:24] = '{
    // Filter 0
    '{
        {16'hACEA, 16'h3678, 16'h33E7, 16'hB606, 16'hB3C7, 16'h22BE, 16'h3529, 16'hA874, 16'hB521, 16'hB28F, 16'hA056, 16'h3406, 16'hA90B, 16'h3112, 16'h2533, 16'h319C, 16'hA1BF, 16'hA105, 16'h2D39, 16'hAC84, 16'h31A1, 16'hA0E6, 16'h9AE1, 16'h30C8, 16'h2E81}
    },
    // Filter 1
    '{
        {16'h31E5, 16'h3542, 16'h36B2, 16'h31F9, 16'hAE40, 16'hB71D, 16'hB5E7, 16'hB4E5, 16'hACCC, 16'h2B28, 16'hB11A, 16'hB611, 16'hB541, 16'hA9FB, 16'h2D56, 16'hB19F, 16'hB25A, 16'h3661, 16'h2C89, 16'hB1C0, 16'h38F3, 16'h38B0, 16'h2E98, 16'hB041, 16'h33B7}
    },
    // Filter 2
    '{
        {16'hAEB9, 16'h2DB0, 16'h2772, 16'hB000, 16'hB055, 16'h31FE, 16'h2FBB, 16'hB590, 16'hB7B0, 16'hAC06, 16'h3334, 16'hB6F8, 16'hB71D, 16'hB422, 16'h341F, 16'hB496, 16'hB826, 16'hB132, 16'h2F9F, 16'h3328, 16'hB439, 16'hB2B7, 16'h2E95, 16'h2CBA, 16'h346C}
    },
    // Filter 3
    '{
        {16'hA973, 16'h33C5, 16'h34F5, 16'h3621, 16'h3675, 16'hAC4C, 16'h36B9, 16'h2FC5, 16'hB3D7, 16'hB0A2, 16'h355A, 16'h312D, 16'hB00E, 16'hB01A, 16'hB466, 16'h3287, 16'hB4F3, 16'hB6F8, 16'hB53D, 16'hB122, 16'hB6B1, 16'hA5DD, 16'h3096, 16'h328D, 16'hAA92}
    }
};

localparam [15:0] BIASES[0:3] = '{16'h2B8C, 16'hB429, 16'hBE68, 16'h2C85};
